// test sv
